module a(
    a,
);
endmodule